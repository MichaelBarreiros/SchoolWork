/*****************************************************************************
 *                                                                           *
 * Module:       Lab5                                                        *
 * Description:                                                              *
 *      This module is the top level module of 2DA4 lab 5                    *
 *                                                                           *
 *****************************************************************************/

module lab5 (
input				CLOCK_50,	
input		[0:0]	KEY, 
input 	[7:0] SW,               //for reset
output 	[7:0] LEDR,

// Bidirectionals
inout		[15:0]	DRAM_DQ,

// Outputs

output		[12:0]	DRAM_ADDR,
output 		[1:0]		DRAM_BA,
output					DRAM_LDQM,  //data mask; when it is low, the DQ is valid for reading and writing. 
output					DRAM_UDQM,
output					DRAM_RAS_N,
output 					DRAM_CAS_N,
output 					DRAM_CLK,
output					DRAM_CKE,
output 					DRAM_WE_N,
output 					DRAM_CS_N


);


// Internal Wires
wire		[12:0]	address;
wire		[1:0]		byte_enable;
wire					rw;
wire		[15:0]	write_data;
wire		[15:0]	read_data;

// The following dummy wires are there just to ensure that 
// Quartus does not perform certain optimizations, which may
// result in these signals appearing inverted when observed in SignalTap II
// The key to this is the /*synthesis keep */ comment, which actually
// has a meaning to Quartus. It is important that the comment appear before the semicolon
// This comment does not affect functionality in any significant way
wire				DRAM_CS_N_wire /*synthesis keep */;
wire				DRAM_WE_N_wire /*synthesis keep */;
wire				DRAM_UDQM_wire /*synthesis keep */;
wire				DRAM_LDQM_wire /*synthesis keep */;


//assign DRAM_CS_N = DRAM_CS_N_wire;
//assign DRAM_WE_N = DRAM_WE_N_wire;
//assign DRAM_UB_N = DRAM_UDQM_wire;
//assign DRAM_LB_N = DRAM_LDQM_wire;

assign LEDR=SW;


//Instantiate your sopc_system module generated by Qsys.  

sopc_system NiosII (
		.clk_clk           (CLOCK_50),           //        clk.clk
		.reset_reset_n     (KEY),     //      reset.reset_n
		.dram_addr_export  (DRAM_ADDR),  //  dram_addr.export
		.dram_ba_export    (DRAM_BA),    //    dram_ba.export
		.dram_cas_n_export (DRAM_CAS_N), // dram_cas_n.export
		.dram_cke_export   (DRAM_CKE),   //   dram_cke.export
		.dram_cs_n_export  (DRAM_CS_N),  //  dram_cs_n.export
		.dram_dq_export    (DRAM_DQ),    //    dram_dq.export
		.dram_ldqm_export  (DRAM_LDQM),  //  dram_ldqm.export
		.dram_ras_n_export (DRAM_RAS_N), // dram_ras_n.export
		.dram_udqm_export  (DRAM_UDQM),  //  dram_udqm.export
		.dram_we_n_export  (DRAM_WE_N),  //  dram_we_n.export
		.sdram_clk_clk     (DRAM_CLK));     //  sdram_clk.clk
endmodule
