module lab1 (x1, x2, x3, x4, f1, f2);
	input x1, x2, x3, x4;
	output f1, f2;
	assign X = x1x2;
	assign Y = y1y2;

		
	assign f1 = (X != Y);
	assign f2 = (X >= Y);
endmodule
